/*
 * user_module_341263346544149074.v
 */

`default_nettype none

module user_module_341263346544149074 (
	input  wire  [7:0] io_in,
	output wire  [7:0] io_out
);

	assign io_out = io_in;

endmodule // user_module_341263346544149074
